module MAC(
input [7:0] A, B,
input  clk, aclr,
output [15:0] MAC_OUT
);
wire [15:0] MUL_OUT;

endmodule
