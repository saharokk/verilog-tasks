module Demux_1_8(Q, Out, Addr, EN
input Q, EN,
input [2:0] Addr,
output [7:0]Out),
);

endmodule;
